`define VERILATOR 1
